library ieee;
use ieee.std_logic_1164.all;

entity bitwise_identity is
	port (
		a : in std_logic_vector(3 downto 0);
		s : out std_logic_vector(3 downto 0)
	);
end bitwise_identity;

architecture behavioral of bitwise_identity is

begin
	
	s <= a;

end architecture behavioral;